`timescale 1ns / 1ps

module instrMem(
    input   [31:0]  iaddr, // Instruction address
    output  reg [31:0]  dout // Data output (instruction)
    output reg [31:0] nextInstr
    );

    wire [29:0] addr; // Reduced address for word-aligned indexing (30 bits for a larger address range)

    assign addr = iaddr[31:2]; // Word-aligned address (ignoring byte offset)

    

    // Combinational logic for ROM
    always @(*) begin
        case (addr)
            30'd0  : dout = 32'b0000000_01010_00000_000_00100_0010011; // ADDI x4, x0, 10
            30'd1  : dout = 32'b0000001_00000_00100_000_11100_1100011; // BEQ x4, x0, Load
            30'd2  : dout = 32'b1111111_11111_00100_000_00100_0010011; // ADDI x4, x4, -1
            30'd3  : dout = 32'b0000001_00100_00000_000_00101_0010011; // ADDI x5, x0, 36
            30'd4  : dout = 32'b1111111_11100_00101_000_00110_0010011; // ADDI x6, x5, -4
            30'd5  : dout = 32'b1111111_00000_00101_000_10001_1100011; // BEQ x5, x0, Sort
            30'd6  : dout = 32'b0000000_00000_00101_010_00111_0000011; // LW x7, 0(x5)
            30'd7  : dout = 32'b0000000_00000_00110_010_01000_0000011; // LW x8, 0(x6)
            30'd8  : dout = 32'b0000000_00111_01000_010_01001_0110011; // SLT x9, x8, x7
            30'd9  : dout = 32'b0000000_00000_01001_001_01100_1100011; // BNE x9, x0, Not Swap
            30'd10 : dout = 32'b0000000_01000_00101_010_00000_0100011; // SW x8, 0(x5)
            30'd11 : dout = 32'b0000000_00111_00110_010_00000_0100011; // SW x7, 0(x6)
            30'd12 : dout = 32'b1111111_11100_00101_000_00101_0010011; // ADDI x5, x5, -4
            30'd13 : dout = 32'b1111111_11100_00101_000_00110_0010011; // ADDI x6, x5, -4
            30'd14 : dout = 32'b1111110_11101_11111_111_01010_1101111; // JAL x10, Itr
            30'd15 : dout = 32'b0000000_00000_00000_010_00001_0000011; // LW x1, 0(x0)
            30'd16 : dout = 32'b0000000_00100_00000_010_00010_0000011; // LW x2, 4(x0)
            30'd17 : dout = 32'b0000000_01000_00000_010_00011_0000011; // LW x3, 8(x0)
            30'd18 : dout = 32'b0000000_01100_00000_010_00100_0000011; // LW x4, 12(x0)
            30'd19 : dout = 32'b0000000_10000_00000_010_00101_0000011; // LW x5, 16(x0)
            30'd20 : dout = 32'b0000000_10100_00000_010_00110_0000011; // LW x6, 20(x0)
            30'd21 : dout = 32'b0000000_11000_00000_010_00111_0000011; // LW x7, 24(x0)
            30'd22 : dout = 32'b0000000_11100_00000_010_01000_0000011; // LW x8, 28(x0)
            30'd23 : dout = 32'b0000001_00000_00000_010_01001_0000011; // LW x9, 32(x0)
            30'd24 : dout = 32'b0000001_00100_00000_010_01010_0000011; // LW x10, 36(x0)
            default: dout = 32'b00000000_00000000_00000000_00000000;  // Default to NOP
        endcase
    end

endmodule
